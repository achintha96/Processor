module IRAM (
input wire [7:0] address,
input clock,
output reg [15:0] q);

reg [15:0] IRAM [4095:0];

initial begin
    IRAM[0] = 16'b1100000011111111;
    IRAM[1] = 16'b0011000100000010;
    IRAM[2] = 16'b1001101000000000;
    IRAM[3] = 16'b1001110000000000;
    IRAM[4] = 16'b1001100100000000;
    IRAM[5] = 16'b1001101100000000;
    IRAM[6] = 16'b0001001000000000;
    IRAM[7] = 16'b0011010100000110;
    IRAM[8] = 16'b1010101000000000;
    IRAM[9] = 16'b0001001000000000;
    IRAM[10] = 16'b0011010100000110;
    IRAM[11] = 16'b1010101000000000;
    IRAM[12] = 16'b0001001000000000;
    IRAM[13] = 16'b0011010100000110;
    IRAM[14] = 16'b0011011100000001;
    IRAM[15] = 16'b0111001000000000;
    IRAM[16] = 16'b0101100000000000;
    IRAM[17] = 16'b0101011000000000;
    IRAM[18] = 16'b1000010000000000;
    IRAM[19] = 16'b1010110000000000;
    IRAM[20] = 16'b0011000100000101;
    IRAM[21] = 16'b0010001000000000;
    IRAM[22] = 16'b0011001000000001;
    IRAM[23] = 16'b0110101000000000;
    IRAM[24] = 16'b0100000100001011;
    IRAM[25] = 16'b1001101000000000;
    IRAM[26] = 16'b1001110000000000;
    IRAM[27] = 16'b0011100100000001;
    IRAM[28] = 16'b0110001000000000;
    IRAM[29] = 16'b0100001000100001;
    IRAM[30] = 16'b1010101100000000;
    IRAM[31] = 16'b1010100100000000;
    IRAM[32] = 16'b0100000000000110;
    IRAM[33] = 16'b0000000000000000;
    IRAM[34] = 16'b1001101000000000;
    IRAM[35] = 16'b1001110000000000;
    IRAM[36] = 16'b1001100100000000;
    IRAM[37] = 16'b1001101100000000;
    IRAM[38] = 16'b0001001000000000;
    IRAM[39] = 16'b0011010100000110;
    IRAM[40] = 16'b1010100100000000;
    IRAM[41] = 16'b0001001000000000;
    IRAM[42] = 16'b0011010100000110;
    IRAM[43] = 16'b1010100100000000;
    IRAM[44] = 16'b0001001000000000;
    IRAM[45] = 16'b0011010100000110;
    IRAM[46] = 16'b0011011100000001;
    IRAM[47] = 16'b0111001000000000;
    IRAM[48] = 16'b0101100000000000;
    IRAM[49] = 16'b0101011000000000;
    IRAM[50] = 16'b1000010000000000;
    IRAM[51] = 16'b1010101100000000;
    IRAM[52] = 16'b0011000100000101;
    IRAM[53] = 16'b0010001000000000;
    IRAM[54] = 16'b0011100100000001;
    IRAM[55] = 16'b0110001000000000;
    IRAM[56] = 16'b0100000100101011;
    IRAM[57] = 16'b1001100100000000;
    IRAM[58] = 16'b1001101100000000;
    IRAM[59] = 16'b0011101000000001;
    IRAM[60] = 16'b0110001000000000;
    IRAM[61] = 16'b0100001001000001;
    IRAM[62] = 16'b1010110000000000;
    IRAM[63] = 16'b1010101000000000;
    IRAM[64] = 16'b0100000000100110;
    IRAM[65] = 16'b0000000000000000;
    IRAM[66] = 16'b1001110000000000;
    IRAM[67] = 16'b1001101100000000;
    IRAM[68] = 16'b1001101000000000;
    IRAM[69] = 16'b1001100100000000;
    IRAM[70] = 16'b1100000000000010;
    IRAM[71] = 16'b0011000100000011;
    IRAM[72] = 16'b1100000011111110;
    IRAM[73] = 16'b0011000100000010;
    IRAM[74] = 16'b0001001000000000;
    IRAM[75] = 16'b0010001000000000;
    IRAM[76] = 16'b0011101000000001;
    IRAM[77] = 16'b0110001000000000;
    IRAM[78] = 16'b1010110000000000;
    IRAM[79] = 16'b0100001001010011;
    IRAM[80] = 16'b1010101000000000;
    IRAM[81] = 16'b1010101000000000;
    IRAM[82] = 16'b0100000001001010;
    IRAM[83] = 16'b1001101000000000;
    IRAM[84] = 16'b1001110000000000;
    IRAM[85] = 16'b1010101100000000;
    IRAM[86] = 16'b0011100100000001;
    IRAM[87] = 16'b0110001000000000;
    IRAM[88] = 16'b0100001001011100;
    IRAM[89] = 16'b1010100100000000;
    IRAM[90] = 16'b1010100100000000;
    IRAM[91] = 16'b0100000001001010;
    IRAM[92] = 16'b1111000000000000;
end
always @(posedge clock)
begin
	q <= IRAM[address];
end
endmodule